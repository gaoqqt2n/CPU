address <= 
    begin
        100 : x"00000000";
        100 : x"00000004";
        100 : x"0000000c";
    end;
    

        